//******************************************************************************
// file header
//******************************************************************************
//
//  File name: clk_gated.v
//
//  Description: clock gated with enable signal
//
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None


//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module clk_gated (
    clk,
    rst_n,

    mode_i,
    en_ip_i,
    en_i,

    clk_gated_o 
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input clk;
input rst_n;

input [1:0] mode_i;
input en_ip_i;
input en_i;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output clk_gated_o;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
wire en_gated_clk;
wire sel_gated; // 1'b0 -> en_ip_i, 1'b1 -> ram enable_singal(en_i)

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg en_clk; // clk enable signal(negedge clk sampled)

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
assign clk_gated_o = en_clk & clk;

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
assign en_gated_clk = mode_i[1];
assign sel_gated = mode_i[0];

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (negedge clk or negedge rst_n) begin
    if (!rst_n)
        en_clk <= #TD 1'b0;
    else if (!en_gated_clk)
             en_clk <= #TD 1'b1;
         else if (sel_gated)
                  en_clk <= #TD en_i;
              else
                  en_clk <= #TD en_ip_i;
end

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
