//******************************************************************************
// file header
//******************************************************************************
//
//  File name: ctrl_sync.v
//
//  Description:
//
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None


//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module ctrl_sync (
    clk_src,
    clk_dest,
    rst_src_n,
    rst_dest_n,

    ctrl_i,

    ctrl_sync_o
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
parameter FAST2SLOW = 0;

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input clk_src;
input clk_dest;
input rst_src_n;
input rst_dest_n;

input ctrl_i;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output ctrl_sync_o;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
wire ctrl_src; // ctrl signal will be synchronized to destination clock

wire ctrl_clr; // clear ctrl_lvl after synchronized to destination clock
wire ctrl_flag;

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
reg ctrl_sync_o;

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg ctrl_lvl; // multi clock cycle ctrl

// clear signal for level control
reg clr_ctrl_q;
reg clr_ctrl_q1;

reg ctrl_sync_q;

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
assign ctrl_src = (FAST2SLOW)? ctrl_lvl: ctrl_i;

assign ctrl_clr = clr_ctrl_q1? 1'b0: ctrl_lvl;
assign ctrl_flag = ctrl_i? 1'b1: ctrl_clr;

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
always @ (negedge rst_dest_n or posedge clk_dest) begin
    if (!rst_dest_n)
        ctrl_sync_o <= #TD 1'b0;
    else
        ctrl_sync_o <= #TD ctrl_sync_q;
end

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (negedge rst_src_n or posedge clk_src) begin
    if (!rst_src_n)
        ctrl_lvl <= #TD 1'b0;
    else
        ctrl_lvl <= #TD ctrl_flag;
end

always @ (negedge rst_src_n or posedge clk_src) begin
    if (!rst_src_n)
        clr_ctrl_q <= #TD 1'b0;
    else
        clr_ctrl_q <= #TD ctrl_sync_o;
end

always @ (negedge rst_src_n or posedge clk_src) begin
    if (!rst_src_n)
        clr_ctrl_q1 <= #TD 1'b0;
    else
        clr_ctrl_q1 <= #TD clr_ctrl_q;
end

always @ (negedge rst_dest_n or posedge clk_dest) begin
    if (!rst_dest_n)
        ctrl_sync_q <= #TD 1'b0;
    else
        ctrl_sync_q <= #TD ctrl_src;
end

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
